`timescale 1ns / 1ps

module iir_wishbone_tb;

    // Parameters
    parameter DATA_WIDTH = 32;
    parameter ADDR_WIDTH = 6;
    parameter CLK_PERIOD = 10; // 100 MHz clock (10 ns period)
    parameter SAMPLE_PERIOD = 20833; // 48 kHz sampling period (20833 ns)

    // Signals
    reg wb_clk_i;
    reg wb_rst_i;
    reg [ADDR_WIDTH-1:0] wb_adr_i;
    reg [DATA_WIDTH-1:0] wb_dat_i;
    wire [DATA_WIDTH-1:0] wb_dat_o;
    reg wb_we_i;
    reg wb_stb_i;
    reg wb_cyc_i;
    wire wb_ack_o;

    // Instantiate the Unit Under Test (UUT)
    iir_wishbone #(
        .DATA_WIDTH(DATA_WIDTH),
        .ADDR_WIDTH(ADDR_WIDTH)
    ) DUT (
        .wb_clk_i(wb_clk_i),
        .wb_rst_i(wb_rst_i),
        .wb_adr_i(wb_adr_i),
        .wb_dat_i(wb_dat_i),
        .wb_dat_o(wb_dat_o),
        .wb_we_i(wb_we_i),
        .wb_stb_i(wb_stb_i),
        .wb_cyc_i(wb_cyc_i),
        .wb_ack_o(wb_ack_o)
    );

    // Clock generation
    initial wb_clk_i = 0;
    always #(CLK_PERIOD/2) wb_clk_i = ~wb_clk_i;

    // Wishbone write task
    task wishbone_write;
        input [ADDR_WIDTH-1:0] addr;
        input [DATA_WIDTH-1:0] data;
        begin
            @(posedge wb_clk_i);
            wb_adr_i = addr;
            wb_dat_i = data;
            wb_we_i = 1;
            wb_stb_i = 1;
            wb_cyc_i = 1;
            @(posedge wb_clk_i);
            while (!wb_ack_o) @(posedge wb_clk_i);
            wb_stb_i = 0;
            wb_cyc_i = 0;
        end
    endtask

    // Wishbone read task
    task wishbone_read;
        input [ADDR_WIDTH-1:0] addr;
        output [DATA_WIDTH-1:0] data;
        begin
            @(posedge wb_clk_i);
            wb_adr_i = addr;
            wb_we_i = 0;
            wb_stb_i = 1;
            wb_cyc_i = 1;
            @(posedge wb_clk_i);
            while (!wb_ack_o) @(posedge wb_clk_i);
            data = wb_dat_o;
            wb_stb_i = 0;
            wb_cyc_i = 0;
        end
    endtask

    // Test procedure
    initial begin
        // Initialize signals
        wb_rst_i = 1;
        wb_adr_i = 0;
        wb_dat_i = 0;
        wb_we_i = 0;
        wb_stb_i = 0;
        wb_cyc_i = 0;

        // Reset
        #10;
        wb_rst_i = 1;
        #20;
        wb_rst_i = 0;
        #10;
        wb_rst_i = 1;

        // Initialize coefficients (from original iir.v)
        wishbone_write(6'h00, 5509);    // b0_s1
        wishbone_write(6'h04, 11019);   // b1_s1
        wishbone_write(6'h08, 5509);    // b2_s1
        wishbone_write(6'h0C, -1998080); // a1_s1
        wishbone_write(6'h10, 971584);  // a2_s1
        wishbone_write(6'h14, 5180);    // b0_s2
        wishbone_write(6'h18, 10360);   // b1_s2
        wishbone_write(6'h1C, 5180);    // b2_s2
        wishbone_write(6'h20, -1878592); // delicios
        wishbone_write(6'h24, 850752);  // a2_s2
        wishbone_write(6'h28, 5007);    // b0_s3
        wishbone_write(6'h2C, 10014);   // b1_s3
        wishbone_write(6'h30, 5007);    // b2_s3
        wishbone_write(6'h34, -1815872); // a1_s3
        wishbone_write(6'h38, 787328);  // a2_s3

        // Apply input samples and read outputs
        wishbone_write(6'h3C, 67); #SAMPLE_PERIOD; // Sample(1)
        wishbone_write(6'h3C, -456); #SAMPLE_PERIOD; // Sample(2)
        wishbone_write(6'h3C, 19); #SAMPLE_PERIOD; // Sample(3)
        wishbone_write(6'h3C, 28); #SAMPLE_PERIOD; // Sample(4)
        wishbone_write(6'h3C, 160); #SAMPLE_PERIOD; // Sample(5)
        wishbone_write(6'h3C, 39); #SAMPLE_PERIOD; // Sample(6)
        wishbone_write(6'h3C, 142); #SAMPLE_PERIOD; // Sample(7)
        wishbone_write(6'h3C, 151); #SAMPLE_PERIOD; // Sample(8)
        wishbone_write(6'h3C, 117); #SAMPLE_PERIOD; // Sample(9)
        wishbone_write(6'h3C, 294); #SAMPLE_PERIOD; // Sample(10)
        wishbone_write(6'h3C, 199); #SAMPLE_PERIOD; // Sample(11)
        wishbone_write(6'h3C, 363); #SAMPLE_PERIOD; // Sample(12)
        wishbone_write(6'h3C, 100); #SAMPLE_PERIOD; // Sample(13)
        wishbone_write(6'h3C, 525); #SAMPLE_PERIOD; // Sample(14)
        wishbone_write(6'h3C, 78); #SAMPLE_PERIOD; // Sample(15)
        wishbone_write(6'h3C, 195); #SAMPLE_PERIOD; // Sample(16)
        wishbone_write(6'h3C, -19); #SAMPLE_PERIOD; // Sample(17)
        wishbone_write(6'h3C, 147); #SAMPLE_PERIOD; // Sample(18)
        wishbone_write(6'h3C, 515); #SAMPLE_PERIOD; // Sample(19)
        wishbone_write(6'h3C, 373); #SAMPLE_PERIOD; // Sample(20)
        wishbone_write(6'h3C, 110); #SAMPLE_PERIOD; // Sample(21)
        wishbone_write(6'h3C, 389); #SAMPLE_PERIOD; // Sample(22)
        wishbone_write(6'h3C, 161); #SAMPLE_PERIOD; // Sample(23)
        wishbone_write(6'h3C, -98); #SAMPLE_PERIOD; // Sample(24)
        wishbone_write(6'h3C, 198); #SAMPLE_PERIOD; // Sample(25)
        wishbone_write(6'h3C, 673); #SAMPLE_PERIOD; // Sample(26)
        wishbone_write(6'h3C, 338); #SAMPLE_PERIOD; // Sample(27)
        wishbone_write(6'h3C, -79); #SAMPLE_PERIOD; // Sample(28)
        wishbone_write(6'h3C, 424); #SAMPLE_PERIOD; // Sample(29)
        wishbone_write(6'h3C, 653); #SAMPLE_PERIOD; // Sample(30)
        wishbone_write(6'h3C, 269); #SAMPLE_PERIOD; // Sample(31)
        wishbone_write(6'h3C, 241); #SAMPLE_PERIOD; // Sample(32)
        wishbone_write(6'h3C, 374); #SAMPLE_PERIOD; // Sample(33)
        wishbone_write(6'h3C, 92); #SAMPLE_PERIOD; // Sample(34)
        wishbone_write(6'h3C, 296); #SAMPLE_PERIOD; // Sample(35)
        wishbone_write(6'h3C, 707); #SAMPLE_PERIOD; // Sample(36)
        wishbone_write(6'h3C, 46); #SAMPLE_PERIOD; // Sample(37)
        wishbone_write(6'h3C, 212); #SAMPLE_PERIOD; // Sample(38)
        wishbone_write(6'h3C, 262); #SAMPLE_PERIOD; // Sample(39)
        wishbone_write(6'h3C, 251); #SAMPLE_PERIOD; // Sample(40)
        wishbone_write(6'h3C, 315); #SAMPLE_PERIOD; // Sample(41)
        wishbone_write(6'h3C, 94); #SAMPLE_PERIOD; // Sample(42)
        wishbone_write(6'h3C, -26); #SAMPLE_PERIOD; // Sample(43)
        wishbone_write(6'h3C, 84); #SAMPLE_PERIOD; // Sample(44)
        wishbone_write(6'h3C, -286); #SAMPLE_PERIOD; // Sample(45)
        wishbone_write(6'h3C, 18); #SAMPLE_PERIOD; // Sample(46)
        wishbone_write(6'h3C, 459); #SAMPLE_PERIOD; // Sample(47)
        wishbone_write(6'h3C, -86); #SAMPLE_PERIOD; // Sample(48)
        wishbone_write(6'h3C, 70); #SAMPLE_PERIOD; // Sample(49)
        wishbone_write(6'h3C, 77); #SAMPLE_PERIOD; // Sample(50)
        wishbone_write(6'h3C, 38); #SAMPLE_PERIOD; // Sample(51)
        wishbone_write(6'h3C, -44); #SAMPLE_PERIOD; // Sample(52)
        wishbone_write(6'h3C, -200); #SAMPLE_PERIOD; // Sample(53)
        wishbone_write(6'h3C, -27); #SAMPLE_PERIOD; // Sample(54)
        wishbone_write(6'h3C, -67); #SAMPLE_PERIOD; // Sample(55)
        wishbone_write(6'h3C, -100); #SAMPLE_PERIOD; // Sample(56)
        wishbone_write(6'h3C, -33); #SAMPLE_PERIOD; // Sample(57)
        wishbone_write(6'h3C, -199); #SAMPLE_PERIOD; // Sample(58)
        wishbone_write(6'h3C, -407); #SAMPLE_PERIOD; // Sample(59)
        wishbone_write(6'h3C, -343); #SAMPLE_PERIOD; // Sample(60)
        wishbone_write(6'h3C, -78); #SAMPLE_PERIOD; // Sample(61)
        wishbone_write(6'h3C, -28); #SAMPLE_PERIOD; // Sample(62)
        wishbone_write(6'h3C, -358); #SAMPLE_PERIOD; // Sample(63)
        wishbone_write(6'h3C, -503); #SAMPLE_PERIOD; // Sample(64)
        wishbone_write(6'h3C, -454); #SAMPLE_PERIOD; // Sample(65)
        wishbone_write(6'h3C, -75); #SAMPLE_PERIOD; // Sample(66)
        wishbone_write(6'h3C, -101); #SAMPLE_PERIOD; // Sample(67)
        wishbone_write(6'h3C, -133); #SAMPLE_PERIOD; // Sample(68)
        wishbone_write(6'h3C, -103); #SAMPLE_PERIOD; // Sample(69)
        wishbone_write(6'h3C, -299); #SAMPLE_PERIOD; // Sample(70)
        wishbone_write(6'h3C, -267); #SAMPLE_PERIOD; // Sample(71)
        wishbone_write(6'h3C, -161); #SAMPLE_PERIOD; // Sample(72)
        wishbone_write(6'h3C, -123); #SAMPLE_PERIOD; // Sample(73)
        wishbone_write(6'h3C, 191); #SAMPLE_PERIOD; // Sample(74)
        wishbone_write(6'h3C, -482); #SAMPLE_PERIOD; // Sample(75)
        wishbone_write(6'h3C, -272); #SAMPLE_PERIOD; // Sample(76)
        wishbone_write(6'h3C, -206); #SAMPLE_PERIOD; // Sample(77)
        wishbone_write(6'h3C, -506); #SAMPLE_PERIOD; // Sample(78)
        wishbone_write(6'h3C, -562); #SAMPLE_PERIOD; // Sample(79)
        wishbone_write(6'h3C, -238); #SAMPLE_PERIOD; // Sample(80)
        wishbone_write(6'h3C, -396); #SAMPLE_PERIOD; // Sample(81)
        wishbone_write(6'h3C, -249); #SAMPLE_PERIOD; // Sample(82)
        wishbone_write(6'h3C, -421); #SAMPLE_PERIOD; // Sample(83)
        wishbone_write(6'h3C, -245); #SAMPLE_PERIOD; // Sample(84)
        wishbone_write(6'h3C, -193); #SAMPLE_PERIOD; // Sample(85)
        wishbone_write(6'h3C, -624); #SAMPLE_PERIOD; // Sample(86)
        wishbone_write(6'h3C, -37); #SAMPLE_PERIOD; // Sample(87)
        wishbone_write(6'h3C, -554); #SAMPLE_PERIOD; // Sample(88)
        wishbone_write(6'h3C, -101); #SAMPLE_PERIOD; // Sample(89)
        wishbone_write(6'h3C, -129); #SAMPLE_PERIOD; // Sample(90)
        wishbone_write(6'h3C, -70); #SAMPLE_PERIOD; // Sample(91)
        wishbone_write(6'h3C, 197); #SAMPLE_PERIOD; // Sample(92)
        wishbone_write(6'h3C, -374); #SAMPLE_PERIOD; // Sample(93)
        wishbone_write(6'h3C, -191); #SAMPLE_PERIOD; // Sample(94)
        wishbone_write(6'h3C, -186); #SAMPLE_PERIOD; // Sample(95)
        wishbone_write(6'h3C, 278); #SAMPLE_PERIOD; // Sample(96)
        wishbone_write(6'h3C, 253); #SAMPLE_PERIOD; // Sample(97)
        wishbone_write(6'h3C, 156); #SAMPLE_PERIOD; // Sample(98)
        wishbone_write(6'h3C, -260); #SAMPLE_PERIOD; // Sample(99)
        wishbone_write(6'h3C, -30); #SAMPLE_PERIOD; // Sample(100)
        wishbone_write(6'h3C, 179); #SAMPLE_PERIOD; // Sample(101)
        wishbone_write(6'h3C, 164); #SAMPLE_PERIOD; // Sample(102)
        wishbone_write(6'h3C, -10); #SAMPLE_PERIOD; // Sample(103)
        wishbone_write(6'h3C, 423); #SAMPLE_PERIOD; // Sample(104)
        wishbone_write(6'h3C, 39); #SAMPLE_PERIOD; // Sample(105)
        wishbone_write(6'h3C, 241); #SAMPLE_PERIOD; // Sample(106)
        wishbone_write(6'h3C, 568); #SAMPLE_PERIOD; // Sample(107)
        wishbone_write(6'h3C, 532); #SAMPLE_PERIOD; // Sample(108)
        wishbone_write(6'h3C, 174); #SAMPLE_PERIOD; // Sample(109)
        wishbone_write(6'h3C, 371); #SAMPLE_PERIOD; // Sample(110)
        wishbone_write(6'h3C, 562); #SAMPLE_PERIOD; // Sample(111)
        wishbone_write(6'h3C, 66); #SAMPLE_PERIOD; // Sample(112)
        wishbone_write(6'h3C, 445); #SAMPLE_PERIOD; // Sample(113)
        wishbone_write(6'h3C, 628); #SAMPLE_PERIOD; // Sample(114)
        wishbone_write(6'h3C, 471); #SAMPLE_PERIOD; // Sample(115)
        wishbone_write(6'h3C, 522); #SAMPLE_PERIOD; // Sample(116)
        wishbone_write(6'h3C, 290); #SAMPLE_PERIOD; // Sample(117)
        wishbone_write(6'h3C, 47); #SAMPLE_PERIOD; // Sample(118)
        wishbone_write(6'h3C, 157); #SAMPLE_PERIOD; // Sample(119)
        wishbone_write(6'h3C, 597); #SAMPLE_PERIOD; // Sample(120)
        wishbone_write(6'h3C, 314); #SAMPLE_PERIOD; // Sample(121)
        wishbone_write(6'h3C, 458); #SAMPLE_PERIOD; // Sample(122)
        wishbone_write(6'h3C, 102); #SAMPLE_PERIOD; // Sample(123)
        wishbone_write(6'h3C, -47); #SAMPLE_PERIOD; // Sample(124)
        wishbone_write(6'h3C, -105); #SAMPLE_PERIOD; // Sample(125)
        wishbone_write(6'h3C, 338); #SAMPLE_PERIOD; // Sample(126)
        wishbone_write(6'h3C, -133); #SAMPLE_PERIOD; // Sample(127)
        wishbone_write(6'h3C, 543); #SAMPLE_PERIOD; // Sample(128)
        wishbone_write(6'h3C, 479); #SAMPLE_PERIOD; // Sample(129)
        wishbone_write(6'h3C, 307); #SAMPLE_PERIOD; // Sample(130)
        wishbone_write(6'h3C, 435); #SAMPLE_PERIOD; // Sample(131)
        wishbone_write(6'h3C, 206); #SAMPLE_PERIOD; // Sample(132)
        wishbone_write(6'h3C, -133); #SAMPLE_PERIOD; // Sample(133)
        wishbone_write(6'h3C, 174); #SAMPLE_PERIOD; // Sample(134)
        wishbone_write(6'h3C, 55); #SAMPLE_PERIOD; // Sample(135)
        wishbone_write(6'h3C, 405); #SAMPLE_PERIOD; // Sample(136)
        wishbone_write(6'h3C, 216); #SAMPLE_PERIOD; // Sample(137)
        wishbone_write(6'h3C, 211); #SAMPLE_PERIOD; // Sample(138)
        wishbone_write(6'h3C, 45); #SAMPLE_PERIOD; // Sample(139)
        wishbone_write(6'h3C, -72); #SAMPLE_PERIOD; // Sample(140)
        wishbone_write(6'h3C, 131); #SAMPLE_PERIOD; // Sample(141)
        wishbone_write(6'h3C, -23); #SAMPLE_PERIOD; // Sample(142)
        wishbone_write(6'h3C, 301); #SAMPLE_PERIOD; // Sample(143)
        wishbone_write(6'h3C, -49); #SAMPLE_PERIOD; // Sample(144)
        wishbone_write(6'h3C, -150); #SAMPLE_PERIOD; // Sample(145)
        wishbone_write(6'h3C, -61); #SAMPLE_PERIOD; // Sample(146)
        wishbone_write(6'h3C, 165); #SAMPLE_PERIOD; // Sample(147)
        wishbone_write(6'h3C, -166); #SAMPLE_PERIOD; // Sample(148)
        wishbone_write(6'h3C, -96); #SAMPLE_PERIOD; // Sample(149)
        wishbone_write(6'h3C, -374); #SAMPLE_PERIOD; // Sample(150)
        wishbone_write(6'h3C, -92); #SAMPLE_PERIOD; // Sample(151)
        wishbone_write(6'h3C, -205); #SAMPLE_PERIOD; // Sample(152)
        wishbone_write(6'h3C, -234); #SAMPLE_PERIOD; // Sample(153)
        wishbone_write(6'h3C, -140); #SAMPLE_PERIOD; // Sample(154)
        wishbone_write(6'h3C, -178); #SAMPLE_PERIOD; // Sample(155)
        wishbone_write(6'h3C, -198); #SAMPLE_PERIOD; // Sample(156)
        wishbone_write(6'h3C, 354); #SAMPLE_PERIOD; // Sample(157)
        wishbone_write(6'h3C, -29); #SAMPLE_PERIOD; // Sample(158)
        wishbone_write(6'h3C, 80); #SAMPLE_PERIOD; // Sample(159)
        wishbone_write(6'h3C, 65); #SAMPLE_PERIOD; // Sample(160)
        wishbone_write(6'h3C, -314); #SAMPLE_PERIOD; // Sample(161)
        wishbone_write(6'h3C, -361); #SAMPLE_PERIOD; // Sample(162)
        wishbone_write(6'h3C, -591); #SAMPLE_PERIOD; // Sample(163)
        wishbone_write(6'h3C, -467); #SAMPLE_PERIOD; // Sample(164)
        wishbone_write(6'h3C, -344); #SAMPLE_PERIOD; // Sample(165)
        wishbone_write(6'h3C, -311); #SAMPLE_PERIOD; // Sample(166)
        wishbone_write(6'h3C, -236); #SAMPLE_PERIOD; // Sample(167)
        wishbone_write(6'h3C, -270); #SAMPLE_PERIOD; // Sample(168)
        wishbone_write(6'h3C, -525); #SAMPLE_PERIOD; // Sample(169)
        wishbone_write(6'h3C, -361); #SAMPLE_PERIOD; // Sample(170)
        wishbone_write(6'h3C, 30); #SAMPLE_PERIOD; // Sample(171)
        wishbone_write(6'h3C, -351); #SAMPLE_PERIOD; // Sample(172)
        wishbone_write(6'h3C, -464); #SAMPLE_PERIOD; // Sample(173)
        wishbone_write(6'h3C, -332); #SAMPLE_PERIOD; // Sample(174)
        wishbone_write(6'h3C, -214); #SAMPLE_PERIOD; // Sample(175)
        wishbone_write(6'h3C, -342); #SAMPLE_PERIOD; // Sample(176)
        wishbone_write(6'h3C, -341); #SAMPLE_PERIOD; // Sample(177)
        wishbone_write(6'h3C, -314); #SAMPLE_PERIOD; // Sample(178)
        wishbone_write(6'h3C, -13); #SAMPLE_PERIOD; // Sample(179)
        wishbone_write(6'h3C, -67); #SAMPLE_PERIOD; // Sample(180)
        wishbone_write(6'h3C, -354); #SAMPLE_PERIOD; // Sample(181)
        wishbone_write(6'h3C, -339); #SAMPLE_PERIOD; // Sample(182)
        wishbone_write(6'h3C, -512); #SAMPLE_PERIOD; // Sample(183)
        wishbone_write(6'h3C, 46); #SAMPLE_PERIOD; // Sample(184)
        wishbone_write(6'h3C, -170); #SAMPLE_PERIOD; // Sample(185)
        wishbone_write(6'h3C, -179); #SAMPLE_PERIOD; // Sample(186)
        wishbone_write(6'h3C, -81); #SAMPLE_PERIOD; // Sample(187)
        wishbone_write(6'h3C, -342); #SAMPLE_PERIOD; // Sample(188)
        wishbone_write(6'h3C, -252); #SAMPLE_PERIOD; // Sample(189)
        wishbone_write(6'h3C, -24); #SAMPLE_PERIOD; // Sample(190)
        wishbone_write(6'h3C, -100); #SAMPLE_PERIOD; // Sample(191)
        wishbone_write(6'h3C, -409); #SAMPLE_PERIOD; // Sample(192)
        wishbone_write(6'h3C, -146); #SAMPLE_PERIOD; // Sample(193)
        wishbone_write(6'h3C, 70); #SAMPLE_PERIOD; // Sample(194)
        wishbone_write(6'h3C, 242); #SAMPLE_PERIOD; // Sample(195)
        wishbone_write(6'h3C, 76); #SAMPLE_PERIOD; // Sample(196)
        wishbone_write(6'h3C, 105); #SAMPLE_PERIOD; // Sample(197)
        wishbone_write(6'h3C, 5); #SAMPLE_PERIOD; // Sample(198)
        wishbone_write(6'h3C, 155); #SAMPLE_PERIOD; // Sample(199)
        wishbone_write(6'h3C, 236); #SAMPLE_PERIOD; // Sample(200)
        wishbone_write(6'h3C, -21); #SAMPLE_PERIOD; // Sample(201)
        wishbone_write(6'h3C, 366); #SAMPLE_PERIOD; // Sample(202)
        wishbone_write(6'h3C, -132); #SAMPLE_PERIOD; // Sample(203)
        wishbone_write(6'h3C, 189); #SAMPLE_PERIOD; // Sample(204)
        wishbone_write(6'h3C, 168); #SAMPLE_PERIOD; // Sample(205)
        wishbone_write(6'h3C, 538); #SAMPLE_PERIOD; // Sample(206)
        wishbone_write(6'h3C, 179); #SAMPLE_PERIOD; // Sample(207)
        wishbone_write(6'h3C, 861); #SAMPLE_PERIOD; // Sample(208)
        wishbone_write(6'h3C, 208); #SAMPLE_PERIOD; // Sample(209)
        wishbone_write(6'h3C, 133); #SAMPLE_PERIOD; // Sample(210)
        wishbone_write(6'h3C, 718); #SAMPLE_PERIOD; // Sample(211)
        wishbone_write(6'h3C, 280); #SAMPLE_PERIOD; // Sample(212)
        wishbone_write(6'h3C, 241); #SAMPLE_PERIOD; // Sample(213)
        wishbone_write(6'h3C, 322); #SAMPLE_PERIOD; // Sample(214)
        wishbone_write(6'h3C, 107); #SAMPLE_PERIOD; // Sample(215)
        wishbone_write(6'h3C, 22); #SAMPLE_PERIOD; // Sample(216)
        wishbone_write(6'h3C, 178); #SAMPLE_PERIOD; // Sample(217)
        wishbone_write(6'h3C, 312); #SAMPLE_PERIOD; // Sample(218)
        wishbone_write(6'h3C, 514); #SAMPLE_PERIOD; // Sample(219)
        wishbone_write(6'h3C, 524); #SAMPLE_PERIOD; // Sample(220)
        wishbone_write(6'h3C, 381); #SAMPLE_PERIOD; // Sample(221)
        wishbone_write(6'h3C, 511); #SAMPLE_PERIOD; // Sample(222)
        wishbone_write(6'h3C, 775); #SAMPLE_PERIOD; // Sample(223)
        wishbone_write(6'h3C, 393); #SAMPLE_PERIOD; // Sample(224)
        wishbone_write(6'h3C, 443); #SAMPLE_PERIOD; // Sample(225)
        wishbone_write(6'h3C, 192); #SAMPLE_PERIOD; // Sample(226)
        wishbone_write(6'h3C, 466); #SAMPLE_PERIOD; // Sample(227)
        wishbone_write(6'h3C, 12); #SAMPLE_PERIOD; // Sample(228)
        wishbone_write(6'h3C, 149); #SAMPLE_PERIOD; // Sample(229)
        wishbone_write(6'h3C, 35); #SAMPLE_PERIOD; // Sample(230)
        wishbone_write(6'h3C, 77); #SAMPLE_PERIOD; // Sample(231)
        wishbone_write(6'h3C, 545); #SAMPLE_PERIOD; // Sample(232)
        wishbone_write(6'h3C, 111); #SAMPLE_PERIOD; // Sample(233)
        wishbone_write(6'h3C, 52); #SAMPLE_PERIOD; // Sample(234)
        wishbone_write(6'h3C, 311); #SAMPLE_PERIOD; // Sample(235)
        wishbone_write(6'h3C, 36); #SAMPLE_PERIOD; // Sample(236)
        wishbone_write(6'h3C, 139); #SAMPLE_PERIOD; // Sample(237)
        wishbone_write(6'h3C, 164); #SAMPLE_PERIOD; // Sample(238)
        wishbone_write(6'h3C, -126); #SAMPLE_PERIOD; // Sample(239)
        wishbone_write(6'h3C, -47); #SAMPLE_PERIOD; // Sample(240)
        wishbone_write(6'h3C, 365); #SAMPLE_PERIOD; // Sample(241)
        wishbone_write(6'h3C, 6); #SAMPLE_PERIOD; // Sample(242)
        wishbone_write(6'h3C, 133); #SAMPLE_PERIOD; // Sample(243)
        wishbone_write(6'h3C, 184); #SAMPLE_PERIOD; // Sample(244)
        wishbone_write(6'h3C, 32); #SAMPLE_PERIOD; // Sample(245)
        wishbone_write(6'h3C, -72); #SAMPLE_PERIOD; // Sample(246)
        wishbone_write(6'h3C, 129); #SAMPLE_PERIOD; // Sample(247)
        wishbone_write(6'h3C, -372); #SAMPLE_PERIOD; // Sample(248)
        wishbone_write(6'h3C, 80); #SAMPLE_PERIOD; // Sample(249)
        wishbone_write(6'h3C, -567); #SAMPLE_PERIOD; // Sample(250)
        wishbone_write(6'h3C, -423); #SAMPLE_PERIOD; // Sample(251)
        wishbone_write(6'h3C, -279); #SAMPLE_PERIOD; // Sample(252)
        wishbone_write(6'h3C, -228); #SAMPLE_PERIOD; // Sample(253)
        wishbone_write(6'h3C, -536); #SAMPLE_PERIOD; // Sample(254)
        wishbone_write(6'h3C, -90); #SAMPLE_PERIOD; // Sample(255)
        wishbone_write(6'h3C, -264); #SAMPLE_PERIOD; // Sample(256)
        wishbone_write(6'h3C, -469); #SAMPLE_PERIOD; // Sample(257)
        wishbone_write(6'h3C, -496); #SAMPLE_PERIOD; // Sample(258)
        wishbone_write(6'h3C, -460); #SAMPLE_PERIOD; // Sample(259)
        wishbone_write(6'h3C, -443); #SAMPLE_PERIOD; // Sample(260)
        wishbone_write(6'h3C, -314); #SAMPLE_PERIOD; // Sample(261)
        wishbone_write(6'h3C, -304); #SAMPLE_PERIOD; // Sample(262)
        wishbone_write(6'h3C, -408); #SAMPLE_PERIOD; // Sample(263)
        wishbone_write(6'h3C, -315); #SAMPLE_PERIOD; // Sample(264)
        wishbone_write(6'h3C, -423); #SAMPLE_PERIOD; // Sample(265)
        wishbone_write(6'h3C, -265); #SAMPLE_PERIOD; // Sample(266)
        wishbone_write(6'h3C, -2); #SAMPLE_PERIOD; // Sample(267)
        wishbone_write(6'h3C, -130); #SAMPLE_PERIOD; // Sample(268)
        wishbone_write(6'h3C, -368); #SAMPLE_PERIOD; // Sample(269)
        wishbone_write(6'h3C, -256); #SAMPLE_PERIOD; // Sample(270)
        wishbone_write(6'h3C, -307); #SAMPLE_PERIOD; // Sample(271)
        wishbone_write(6'h3C, -350); #SAMPLE_PERIOD; // Sample(272)
        wishbone_write(6'h3C, -320); #SAMPLE_PERIOD; // Sample(273)
        wishbone_write(6'h3C, -38); #SAMPLE_PERIOD; // Sample(274)
        wishbone_write(6'h3C, -342); #SAMPLE_PERIOD; // Sample(275)
        wishbone_write(6'h3C, -190); #SAMPLE_PERIOD; // Sample(276)
        wishbone_write(6'h3C, -95); #SAMPLE_PERIOD; // Sample(277)
        wishbone_write(6'h3C, -395); #SAMPLE_PERIOD; // Sample(278)
        wishbone_write(6'h3C, -470); #SAMPLE_PERIOD; // Sample(279)
        wishbone_write(6'h3C, -21); #SAMPLE_PERIOD; // Sample(280)
        wishbone_write(6'h3C, -77); #SAMPLE_PERIOD; // Sample(281)
        wishbone_write(6'h3C, -235); #SAMPLE_PERIOD; // Sample(282)
        wishbone_write(6'h3C, 100); #SAMPLE_PERIOD; // Sample(283)
        wishbone_write(6'h3C, -36); #SAMPLE_PERIOD; // Sample(284)
        wishbone_write(6'h3C, -155); #SAMPLE_PERIOD; // Sample(285)
        wishbone_write(6'h3C, -143); #SAMPLE_PERIOD; // Sample(286)
        wishbone_write(6'h3C, -134); #SAMPLE_PERIOD; // Sample(287)
        wishbone_write(6'h3C, -228); #SAMPLE_PERIOD; // Sample(288)
        wishbone_write(6'h3C, 519); #SAMPLE_PERIOD; // Sample(289)
        wishbone_write(6'h3C, -412); #SAMPLE_PERIOD; // Sample(290)
        wishbone_write(6'h3C, 91); #SAMPLE_PERIOD; // Sample(291)
        wishbone_write(6'h3C, 60); #SAMPLE_PERIOD; // Sample(292)
        wishbone_write(6'h3C, -166); #SAMPLE_PERIOD; // Sample(293)
        wishbone_write(6'h3C, 68); #SAMPLE_PERIOD; // Sample(294)
        wishbone_write(6'h3C, 189); #SAMPLE_PERIOD; // Sample(295)
        wishbone_write(6'h3C, 328); #SAMPLE_PERIOD; // Sample(296)
        wishbone_write(6'h3C, 171); #SAMPLE_PERIOD; // Sample(297)
        wishbone_write(6'h3C, 278); #SAMPLE_PERIOD; // Sample(298)
        wishbone_write(6'h3C, 516); #SAMPLE_PERIOD; // Sample(299)
        wishbone_write(6'h3C, 177); #SAMPLE_PERIOD; // Sample(300)
        wishbone_write(6'h3C, 103); #SAMPLE_PERIOD; // Sample(301)
        wishbone_write(6'h3C, -46); #SAMPLE_PERIOD; // Sample(302)
        wishbone_write(6'h3C, 399); #SAMPLE_PERIOD; // Sample(303)
        wishbone_write(6'h3C, 152); #SAMPLE_PERIOD; // Sample(304)
        wishbone_write(6'h3C, 530); #SAMPLE_PERIOD; // Sample(305)
        wishbone_write(6'h3C, 283); #SAMPLE_PERIOD; // Sample(306)
        wishbone_write(6'h3C, 251); #SAMPLE_PERIOD; // Sample(307)
        wishbone_write(6'h3C, 177); #SAMPLE_PERIOD; // Sample(308)
        wishbone_write(6'h3C, 192); #SAMPLE_PERIOD; // Sample(309)
        wishbone_write(6'h3C, 54); #SAMPLE_PERIOD; // Sample(310)
        wishbone_write(6'h3C, 411); #SAMPLE_PERIOD; // Sample(311)
        wishbone_write(6'h3C, 219); #SAMPLE_PERIOD; // Sample(312)
        wishbone_write(6'h3C, 421); #SAMPLE_PERIOD; // Sample(313)
        wishbone_write(6'h3C, -22); #SAMPLE_PERIOD; // Sample(314)
        wishbone_write(6'h3C, 362); #SAMPLE_PERIOD; // Sample(315)
        wishbone_write(6'h3C, 120); #SAMPLE_PERIOD; // Sample(316)
        wishbone_write(6'h3C, -7); #SAMPLE_PERIOD; // Sample(317)
        wishbone_write(6'h3C, 239); #SAMPLE_PERIOD; // Sample(318)
        wishbone_write(6'h3C, 394); #SAMPLE_PERIOD; // Sample(319)
        wishbone_write(6'h3C, 465); #SAMPLE_PERIOD; // Sample(320)
        wishbone_write(6'h3C, 494); #SAMPLE_PERIOD; // Sample(321)
        wishbone_write(6'h3C, 177); #SAMPLE_PERIOD; // Sample(322)
        wishbone_write(6'h3C, 56); #SAMPLE_PERIOD; // Sample(323)
        wishbone_write(6'h3C, 802); #SAMPLE_PERIOD; // Sample(324)
        wishbone_write(6'h3C, 108); #SAMPLE_PERIOD; // Sample(325)
        wishbone_write(6'h3C, 64); #SAMPLE_PERIOD; // Sample(326)
        wishbone_write(6'h3C, 273); #SAMPLE_PERIOD; // Sample(327)
        wishbone_write(6'h3C, -37); #SAMPLE_PERIOD; // Sample(328)
        wishbone_write(6'h3C, 24); #SAMPLE_PERIOD; // Sample(329)
        wishbone_write(6'h3C, -156); #SAMPLE_PERIOD; // Sample(330)
        wishbone_write(6'h3C, 77); #SAMPLE_PERIOD; // Sample(331)
        wishbone_write(6'h3C, -117); #SAMPLE_PERIOD; // Sample(332)
        wishbone_write(6'h3C, 152); #SAMPLE_PERIOD; // Sample(333)
        wishbone_write(6'h3C, 95); #SAMPLE_PERIOD; // Sample(334)
        wishbone_write(6'h3C, -97); #SAMPLE_PERIOD; // Sample(335)
        wishbone_write(6'h3C, -53); #SAMPLE_PERIOD; // Sample(336)
        wishbone_write(6'h3C, -108); #SAMPLE_PERIOD; // Sample(337)
        wishbone_write(6'h3C, 12); #SAMPLE_PERIOD; // Sample(338)
        wishbone_write(6'h3C, -163); #SAMPLE_PERIOD; // Sample(339)
        wishbone_write(6'h3C, -8); #SAMPLE_PERIOD; // Sample(340)
        wishbone_write(6'h3C, -239); #SAMPLE_PERIOD; // Sample(341)
        wishbone_write(6'h3C, 15); #SAMPLE_PERIOD; // Sample(342)
        wishbone_write(6'h3C, -146); #SAMPLE_PERIOD; // Sample(343)
        wishbone_write(6'h3C, -521); #SAMPLE_PERIOD; // Sample(344)
        wishbone_write(6'h3C, -114); #SAMPLE_PERIOD; // Sample(345)
        wishbone_write(6'h3C, 12); #SAMPLE_PERIOD; // Sample(346)
        wishbone_write(6'h3C, 56); #SAMPLE_PERIOD; // Sample(347)
        wishbone_write(6'h3C, -155); #SAMPLE_PERIOD; // Sample(348)
        wishbone_write(6'h3C, 68); #SAMPLE_PERIOD; // Sample(349)
        wishbone_write(6'h3C, -95); #SAMPLE_PERIOD; // Sample(350)
        wishbone_write(6'h3C, 160); #SAMPLE_PERIOD; // Sample(351)
        wishbone_write(6'h3C, -199); #SAMPLE_PERIOD; // Sample(352)
        wishbone_write(6'h3C, -169); #SAMPLE_PERIOD; // Sample(353)
        wishbone_write(6'h3C, -187); #SAMPLE_PERIOD; // Sample(354)
        wishbone_write(6'h3C, -172); #SAMPLE_PERIOD; // Sample(355)
        wishbone_write(6'h3C, -127); #SAMPLE_PERIOD; // Sample(356)
        wishbone_write(6'h3C, -89); #SAMPLE_PERIOD; // Sample(357)
        wishbone_write(6'h3C, -480); #SAMPLE_PERIOD; // Sample(358)
        wishbone_write(6'h3C, -542); #SAMPLE_PERIOD; // Sample(359)
        wishbone_write(6'h3C, -47); #SAMPLE_PERIOD; // Sample(360)
        wishbone_write(6'h3C, -117); #SAMPLE_PERIOD; // Sample(361)
        wishbone_write(6'h3C, -459); #SAMPLE_PERIOD; // Sample(362)
        wishbone_write(6'h3C, -306); #SAMPLE_PERIOD; // Sample(363)
        wishbone_write(6'h3C, 55); #SAMPLE_PERIOD; // Sample(364)
        wishbone_write(6'h3C, -508); #SAMPLE_PERIOD; // Sample(365)
        wishbone_write(6'h3C, -222); #SAMPLE_PERIOD; // Sample(366)
        wishbone_write(6'h3C, -539); #SAMPLE_PERIOD; // Sample(367)
        wishbone_write(6'h3C, -236); #SAMPLE_PERIOD; // Sample(368)
        wishbone_write(6'h3C, -202); #SAMPLE_PERIOD; // Sample(369)
        wishbone_write(6'h3C, -283); #SAMPLE_PERIOD; // Sample(370)
        wishbone_write(6'h3C, -60); #SAMPLE_PERIOD; // Sample(371)
        wishbone_write(6'h3C, -252); #SAMPLE_PERIOD; // Sample(372)
        wishbone_write(6'h3C, 12); #SAMPLE_PERIOD; // Sample(373)
        wishbone_write(6'h3C, 9); #SAMPLE_PERIOD; // Sample(374)
        wishbone_write(6'h3C, -235); #SAMPLE_PERIOD; // Sample(375)
        wishbone_write(6'h3C, -118); #SAMPLE_PERIOD; // Sample(376)
        wishbone_write(6'h3C, -110); #SAMPLE_PERIOD; // Sample(377)
        wishbone_write(6'h3C, 50); #SAMPLE_PERIOD; // Sample(378)
        wishbone_write(6'h3C, 120); #SAMPLE_PERIOD; // Sample(379)
        wishbone_write(6'h3C, 54); #SAMPLE_PERIOD; // Sample(380)
        wishbone_write(6'h3C, -73); #SAMPLE_PERIOD; // Sample(381)
        wishbone_write(6'h3C, -227); #SAMPLE_PERIOD; // Sample(382)
        wishbone_write(6'h3C, -282); #SAMPLE_PERIOD; // Sample(383)
        wishbone_write(6'h3C, 188); #SAMPLE_PERIOD; // Sample(384)
        wishbone_write(6'h3C, 377); #SAMPLE_PERIOD; // Sample(385)
        wishbone_write(6'h3C, 71); #SAMPLE_PERIOD; // Sample(386)
        wishbone_write(6'h3C, 26); #SAMPLE_PERIOD; // Sample(387)
        wishbone_write(6'h3C, 236); #SAMPLE_PERIOD; // Sample(388)
        wishbone_write(6'h3C, -239); #SAMPLE_PERIOD; // Sample(389)
        wishbone_write(6'h3C, 47); #SAMPLE_PERIOD; // Sample(390)
        wishbone_write(6'h3C, -262); #SAMPLE_PERIOD; // Sample(391)
        wishbone_write(6'h3C, 214); #SAMPLE_PERIOD; // Sample(392)
        wishbone_write(6'h3C, 156); #SAMPLE_PERIOD; // Sample(393)
        wishbone_write(6'h3C, 229); #SAMPLE_PERIOD; // Sample(394)
        wishbone_write(6'h3C, 102); #SAMPLE_PERIOD; // Sample(395)
        wishbone_write(6'h3C, -154); #SAMPLE_PERIOD; // Sample(396)
        wishbone_write(6'h3C, 400); #SAMPLE_PERIOD; // Sample(397)
        wishbone_write(6'h3C, 103); #SAMPLE_PERIOD; // Sample(398)
        wishbone_write(6'h3C, 272); #SAMPLE_PERIOD; // Sample(399)
        wishbone_write(6'h3C, 429); #SAMPLE_PERIOD; // Sample(400)
        wishbone_write(6'h3C, 368); #SAMPLE_PERIOD; // Sample(401)
        wishbone_write(6'h3C, 113); #SAMPLE_PERIOD; // Sample(402)
        wishbone_write(6'h3C, 228); #SAMPLE_PERIOD; // Sample(403)
        wishbone_write(6'h3C, 243); #SAMPLE_PERIOD; // Sample(404)
        wishbone_write(6'h3C, 477); #SAMPLE_PERIOD; // Sample(405)
        wishbone_write(6'h3C, 537); #SAMPLE_PERIOD; // Sample(406)
        wishbone_write(6'h3C, 97); #SAMPLE_PERIOD; // Sample(407)
        wishbone_write(6'h3C, 107); #SAMPLE_PERIOD; // Sample(408)
        wishbone_write(6'h3C, 325); #SAMPLE_PERIOD; // Sample(409)
        wishbone_write(6'h3C, 299); #SAMPLE_PERIOD; // Sample(410)
        wishbone_write(6'h3C, 335); #SAMPLE_PERIOD; // Sample(411)
        wishbone_write(6'h3C, 96); #SAMPLE_PERIOD; // Sample(412)
        wishbone_write(6'h3C, 37); #SAMPLE_PERIOD; // Sample(413)
        wishbone_write(6'h3C, 269); #SAMPLE_PERIOD; // Sample(414)
        wishbone_write(6'h3C, 511); #SAMPLE_PERIOD; // Sample(415)
        wishbone_write(6'h3C, 389); #SAMPLE_PERIOD; // Sample(416)
        wishbone_write(6'h3C, 238); #SAMPLE_PERIOD; // Sample(417)
        wishbone_write(6'h3C, 177); #SAMPLE_PERIOD; // Sample(418)
        wishbone_write(6'h3C, 26); #SAMPLE_PERIOD; // Sample(419)
        wishbone_write(6'h3C, 396); #SAMPLE_PERIOD; // Sample(420)
        wishbone_write(6'h3C, 374); #SAMPLE_PERIOD; // Sample(421)
        wishbone_write(6'h3C, 167); #SAMPLE_PERIOD; // Sample(422)
        wishbone_write(6'h3C, 256); #SAMPLE_PERIOD; // Sample(423)
        wishbone_write(6'h3C, 219); #SAMPLE_PERIOD; // Sample(424)
        wishbone_write(6'h3C, 325); #SAMPLE_PERIOD; // Sample(425)
        wishbone_write(6'h3C, 443); #SAMPLE_PERIOD; // Sample(426)
        wishbone_write(6'h3C, -217); #SAMPLE_PERIOD; // Sample(427)
        wishbone_write(6'h3C, 38); #SAMPLE_PERIOD; // Sample(428)
        wishbone_write(6'h3C, 63); #SAMPLE_PERIOD; // Sample(429)
        wishbone_write(6'h3C, -182); #SAMPLE_PERIOD; // Sample(430)
        wishbone_write(6'h3C, -16); #SAMPLE_PERIOD; // Sample(431)
        wishbone_write(6'h3C, 174); #SAMPLE_PERIOD; // Sample(432)
        wishbone_write(6'h3C, -143); #SAMPLE_PERIOD; // Sample(433)
        wishbone_write(6'h3C, -417); #SAMPLE_PERIOD; // Sample(434)
        wishbone_write(6'h3C, -232); #SAMPLE_PERIOD; // Sample(435)
        wishbone_write(6'h3C, -5); #SAMPLE_PERIOD; // Sample(436)
        wishbone_write(6'h3C, -222); #SAMPLE_PERIOD; // Sample(437)
        wishbone_write(6'h3C, 83); #SAMPLE_PERIOD; // Sample(438)
        wishbone_write(6'h3C, -220); #SAMPLE_PERIOD; // Sample(439)
        wishbone_write(6'h3C, -89); #SAMPLE_PERIOD; // Sample(440)
        wishbone_write(6'h3C, -263); #SAMPLE_PERIOD; // Sample(441)
        wishbone_write(6'h3C, -48); #SAMPLE_PERIOD; // Sample(442)
        wishbone_write(6'h3C, -493); #SAMPLE_PERIOD; // Sample(443)
        wishbone_write(6'h3C, 112); #SAMPLE_PERIOD; // Sample(444)
        wishbone_write(6'h3C, -253); #SAMPLE_PERIOD; // Sample(445)
        wishbone_write(6'h3C, -252); #SAMPLE_PERIOD; // Sample(446)
        wishbone_write(6'h3C, -507); #SAMPLE_PERIOD; // Sample(447)
        wishbone_write(6'h3C, -249); #SAMPLE_PERIOD; // Sample(448)
        wishbone_write(6'h3C, -273); #SAMPLE_PERIOD; // Sample(449)
        wishbone_write(6'h3C, -497); #SAMPLE_PERIOD; // Sample(450)
        wishbone_write(6'h3C, -164); #SAMPLE_PERIOD; // Sample(451)
        wishbone_write(6'h3C, 96); #SAMPLE_PERIOD; // Sample(452)
        wishbone_write(6'h3C, -65); #SAMPLE_PERIOD; // Sample(453)
        wishbone_write(6'h3C, -306); #SAMPLE_PERIOD; // Sample(454)
        wishbone_write(6'h3C, -192); #SAMPLE_PERIOD; // Sample(455)
        wishbone_write(6'h3C, -259); #SAMPLE_PERIOD; // Sample(456)
        wishbone_write(6'h3C, -221); #SAMPLE_PERIOD; // Sample(457)
        wishbone_write(6'h3C, -689); #SAMPLE_PERIOD; // Sample(458)
        wishbone_write(6'h3C, -468); #SAMPLE_PERIOD; // Sample(459)
        wishbone_write(6'h3C, -348); #SAMPLE_PERIOD; // Sample(460)
        wishbone_write(6'h3C, -170); #SAMPLE_PERIOD; // Sample(461)
        wishbone_write(6'h3C, -215); #SAMPLE_PERIOD; // Sample(462)
        wishbone_write(6'h3C, -296); #SAMPLE_PERIOD; // Sample(463)
        wishbone_write(6'h3C, -677); #SAMPLE_PERIOD; // Sample(464)
        wishbone_write(6'h3C, -529); #SAMPLE_PERIOD; // Sample(465)
        wishbone_write(6'h3C, 4); #SAMPLE_PERIOD; // Sample(466)
        wishbone_write(6'h3C, -212); #SAMPLE_PERIOD; // Sample(467)
        wishbone_write(6'h3C, -223); #SAMPLE_PERIOD; // Sample(468)
        wishbone_write(6'h3C, -276); #SAMPLE_PERIOD; // Sample(469)
        wishbone_write(6'h3C, 351); #SAMPLE_PERIOD; // Sample(470)
        wishbone_write(6'h3C, -312); #SAMPLE_PERIOD; // Sample(471)
        wishbone_write(6'h3C, -194); #SAMPLE_PERIOD; // Sample(472)
        wishbone_write(6'h3C, -49); #SAMPLE_PERIOD; // Sample(473)
        wishbone_write(6'h3C, 117); #SAMPLE_PERIOD; // Sample(474)
        wishbone_write(6'h3C, -140); #SAMPLE_PERIOD; // Sample(475)
        wishbone_write(6'h3C, 87); #SAMPLE_PERIOD; // Sample(476)
        wishbone_write(6'h3C, 110); #SAMPLE_PERIOD; // Sample(477)
        wishbone_write(6'h3C, -10); #SAMPLE_PERIOD; // Sample(478)
        wishbone_write(6'h3C, -287); #SAMPLE_PERIOD; // Sample(479)
        wishbone_write(6'h3C, 132); #SAMPLE_PERIOD; // Sample(480)
        wishbone_write(6'h3C, 20); #SAMPLE_PERIOD; // Sample(481)
        wishbone_write(6'h3C, 313); #SAMPLE_PERIOD; // Sample(482)
        wishbone_write(6'h3C, -119); #SAMPLE_PERIOD; // Sample(483)
        wishbone_write(6'h3C, 58); #SAMPLE_PERIOD; // Sample(484)
        wishbone_write(6'h3C, -17); #SAMPLE_PERIOD; // Sample(485)
        wishbone_write(6'h3C, -251); #SAMPLE_PERIOD; // Sample(486)
        wishbone_write(6'h3C, -83); #SAMPLE_PERIOD; // Sample(487)
        wishbone_write(6'h3C, -236); #SAMPLE_PERIOD; // Sample(488)
        wishbone_write(6'h3C, 469); #SAMPLE_PERIOD; // Sample(489)
        wishbone_write(6'h3C, 213); #SAMPLE_PERIOD; // Sample(490)
        wishbone_write(6'h3C, 296); #SAMPLE_PERIOD; // Sample(491)
        wishbone_write(6'h3C, 237); #SAMPLE_PERIOD; // Sample(492)
        wishbone_write(6'h3C, 423); #SAMPLE_PERIOD; // Sample(493)
        wishbone_write(6'h3C, 512); #SAMPLE_PERIOD; // Sample(494)
        wishbone_write(6'h3C, 162); #SAMPLE_PERIOD; // Sample(495)
        wishbone_write(6'h3C, 67); #SAMPLE_PERIOD; // Sample(496)
        wishbone_write(6'h3C, 469); #SAMPLE_PERIOD; // Sample(497)
        wishbone_write(6'h3C, 693); #SAMPLE_PERIOD; // Sample(498)
        wishbone_write(6'h3C, 236); #SAMPLE_PERIOD; // Sample(499)
        wishbone_write(6'h3C, 141); #SAMPLE_PERIOD; // Sample(500)

        // Stop simulation
        $stop;
    end

    // Monitor outputs
    reg [DATA_WIDTH-1:0] y_out;
    always @(posedge wb_clk_i) begin
        if (wb_ack_o && !wb_we_i && wb_adr_i == 6'h40) begin
            $display("Time: %0t ns, Output y: %0d", $time, wb_dat_o);
        end
    end

endmodule